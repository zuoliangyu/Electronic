library verilog;
use verilog.vl_types.all;
entity CNT32_vlg_vec_tst is
end CNT32_vlg_vec_tst;
