LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY STM32_OUT1 IS
	GENERIC (ADDR8:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0008";
	ADDR9:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0009");
	PORT(CS,RD,FLAG: IN STD_LOGIC;
	AD_FIFO_DATA:IN STD_LOGIC_VECTOR(13 downto 0);
	ADDR:IN STD_LOGIC_VECTOR(15 downto 0);
	DB:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE BHV OF STM32_OUT1 IS
	
BEGIN
	PROCESS(CS,RD,FLAG,ADDR,AD_FIFO_DATA)
	BEGIN
		IF CS='0' AND RD='0' THEN
				CASE(ADDR) IS
					WHEN ADDR9 => IF FLAG='1' THEN DB<=X"0001";
										ELSE DB<=X"0000"; END IF;
					WHEN ADDR8 => DB<="00" & AD_FIFO_DATA;
					WHEN OTHERS => DB<=(OTHERS=>'Z');
				END CASE;
		ELSE DB<=(OTHERS=>'Z');
		END IF;
	END PROCESS;
END BHV;