--关于接收DSP控制
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
ENTITY DSP_IN IS
	GENERIC (ADDR1:STD_LOGIC_VECTOR(11 DOWNTO 0):=X"001");
	PORT(CS,WR: IN STD_LOGIC;
	DB:IN STD_LOGIC_VECTOR(15 downto 0);
	ADDR:IN STD_LOGIC_VECTOR(11 downto 0);
	DBOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE BHV OF DSP_IN IS
	--SIGNAL Q1,Q1BASE:STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
	PROCESS(CS,WR,ADDR,DB)
	BEGIN
		IF CS='0' AND WR='0' THEN
			IF ADDR=ADDR1 THEN
					DBOUT<=DB;
			END IF;
		END IF;
	END PROCESS;
END BHV;