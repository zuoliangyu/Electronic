LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DS_P_OUT IS
	GENERIC (ADDR2:STD_LOGIC_VECTOR(11 DOWNTO 0):=x"002";
	ADDR3:STD_LOGIC_VECTOR(11 DOWNTO 0):=x"003";
	ADDR4:STD_LOGIC_VECTOR(11 DOWNTO 0):=x"004";
	ADDR5:STD_LOGIC_VECTOR(11 DOWNTO 0):=x"005");
	PORT(CS,WR: IN STD_LOGIC;
	DATA1,DATA2:IN STD_LOGIC_VECTOR(31 downto 0);
	--DATA2:IN STD_LOGIC_VECTOR(31 downto 0);
	ADDR:IN STD_LOGIC_VECTOR(11 downto 0);
	DATAOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE BHV OF DS_P_OUT IS
	
BEGIN
	PROCESS(CS,WR,ADDR,DATA1,DATA2)
	BEGIN
		IF CS='0' THEN
			IF WR='0' THEN
				CASE(ADDR) IS
					WHEN ADDR2 => DATAOUT<=DATA1(31 DOWNTO 16);
					WHEN ADDR3 => DATAOUT<=DATA1(15 DOWNTO 0);
					WHEN ADDR4 => DATAOUT<=DATA2(31 DOWNTO 16);
					WHEN ADDR5 => DATAOUT<=DATA2(15 DOWNTO 0);
					WHEN OTHERS => DATAOUT<=(OTHERS=>'Z');
				END CASE;
			END IF;
		END IF;
	END PROCESS;
END BHV;