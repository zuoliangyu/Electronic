LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY FREQ_DEV IS 
PORT(CLK,EN: IN STD_LOGIC; --输入时钟信号
		FREQH_W,FREQL_W: IN STD_LOGIC_VECTOR(15 DOWNTO 0); -- 频率字
		FREQ_OUT: OUT STD_LOGIC); --分频信号输出
END FREQ_DEV;
ARCHITECTURE DEMO OF FREQ_DEV IS 
	SIGNAL FREQ_WORD: STD_LOGIC_VECTOR(31 DOWNTO 0); 
	SIGNAL ACC:STD_LOGIC_VECTOR(31 DOWNTO 0):=(OTHERS=>'0'); --累加器
	BEGIN 
	PA:PROCESS(CLK,EN,ACC) 
	BEGIN 
		IF(CLK'EVENT AND CLK='1') THEN 
			ACC<=ACC+FREQ_WORD; --累加分频
		END IF; 
		FREQ_OUT<=ACC(31); --最高位输出
	END PROCESS; 
	PB:PROCESS(CLK) --输入频率字的同步化
	BEGIN 
		IF CLK'EVENT AND CLK='1' THEN
			FREQ_WORD<=FREQH_W & FREQL_W;
		END IF;
	END PROCESS;
END DEMO;