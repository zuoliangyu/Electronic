LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
ENTITY CNT32 IS
	PORT(CLR,CLK,CLKBASE,CLKEN,CLKBASEEN: IN STD_LOGIC;
	Q,QBASE:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE BHV OF CNT32 IS
	--SIGNAL Q1,Q1BASE:STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
	A:PROCESS(CLR,CLK,CLKEN)	
	VARIABLE Q1:STD_LOGIC_VECTOR(31 DOWNTO 0);
	BEGIN
	IF CLR='0' THEN Q1:=(OTHERS=>'0');
	ELSIF (CLK'EVENT AND CLK='1') AND CLKEN='1' THEN
		Q1:=Q1+1;
	END IF;	Q<=Q1;
	END PROCESS A;
	B:PROCESS(CLR,CLKBASE,CLKBASEEN)	
	VARIABLE Q1BASE:STD_LOGIC_VECTOR(31 DOWNTO 0);
	BEGIN
	IF CLR='0' THEN  Q1BASE:=(OTHERS=>'0');
	ELSIF (CLKBASE'EVENT AND CLKBASE='1') AND CLKBASEEN='1' THEN	
		Q1BASE:=Q1BASE+1;
	END IF;	QBASE<=Q1BASE;
	END PROCESS B;
END BHV;