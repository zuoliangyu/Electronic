--AD_DIRECT直接采样
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
entity STM32_OUT3 is
	generic (ADDRc:std_logic_vector(15 downto 0):=x"000c";
				ADDRd:std_logic_vector(15 downto 0):=x"000d");
	port(CS,RD,FLAG3 :in std_logic;
			ADDR :in std_logic_vector(15 downto 0);
			DB :out std_logic_vector(15 downto 0);
			AD_FIFO_DATA3 :in std_logic_vector(13 downto 0));
end;
architecture demo of STM32_OUT3 is
begin
	process(CS,RD,ADDR,FLAG3,AD_FIFO_DATA3)
	begin
		if CS='0' and RD='0' then
			case ADDR is
				when ADDRd=> if FLAG3='1' then DB<=x"0001";
								 else DB<=x"0000";end if;
				when ADDRc=> DB<="00" & AD_FIFO_DATA3;
				when others=> DB<="ZZZZZZZZZZZZZZZZ";
			end case;
		else DB<="ZZZZZZZZZZZZZZZZ";
		end if;
	end process;
end demo;