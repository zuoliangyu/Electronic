LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_SIGNED.ALL;
ENTITY STM32_IN IS
	GENERIC (ADDR1:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0001");
	PORT(CS,WR: IN STD_LOGIC;
	DB:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	ADDR:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	DBOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE BHV OF STM32_IN IS
BEGIN
	PROCESS(CS,WR,ADDR,DB)
	BEGIN
		IF CS='0' AND WR='0' THEN
			IF ADDR=ADDR1 THEN
					DBOUT<=DB;
			END IF;
		END IF;
	END PROCESS;
END BHV;