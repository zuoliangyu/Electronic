LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DSP_OUT IS
	GENERIC (ADDR2:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0002";
	ADDR3:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0003";
	ADDR4:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0004";
	ADDR5:STD_LOGIC_VECTOR(15 DOWNTO 0):=x"0005");
	PORT(CS,RD: IN STD_LOGIC;
	DATA1,DATA2:IN STD_LOGIC_VECTOR(31 downto 0);
	ADDR:IN STD_LOGIC_VECTOR(15 downto 0);
	DATAOUT:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END ENTITY;
ARCHITECTURE BHV OF DSP_OUT IS
	
BEGIN
	PROCESS(CS,RD,ADDR,DATA1,DATA2)
	BEGIN
		IF CS='0' AND RD='0' THEN
				CASE(ADDR) IS
					WHEN ADDR2 => DATAOUT<=DATA1(31 DOWNTO 16);
					WHEN ADDR3 => DATAOUT<=DATA1(15 DOWNTO 0);
					WHEN ADDR4 => DATAOUT<=DATA2(31 DOWNTO 16);
					WHEN ADDR5 => DATAOUT<=DATA2(15 DOWNTO 0);
					WHEN OTHERS => DATAOUT<=(OTHERS=>'Z');
				END CASE;
		ELSE DATAOUT<=(OTHERS=>'Z');
		END IF;
	END PROCESS;
END BHV;